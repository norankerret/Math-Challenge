module lab2(x, out);
input [3:0] x;
output [6:0] out;
assign out[0] = ~x[3]&~x[2]&~x[1]&x[0] | ~x[3]&x[2]&~x[1]&~x[0] | x[3]&~x[2]&x[1]&x[0] |
x[3]&x[2]&~x[1]&x[0];
assign out[1] = ~x[3]&x[2]&~x[1]&x[0] | ~x[3]&x[2]&x[1]& ~x[0] | x[3]&~x[2]&x[1]&x[0] |
x[3]&x[2]&~x[1]&~x[0] | x[3]&x[2]&x[1]&~x[0] | x[3]&x[2]&x[1]&x[0];
assign out[2] = ~x[3]&~x[2]&x[1]&~x[0] | x[3]&x[2]&~x[1]&~x[0] | x[3]&x[2]&x[1]&~x[0] |
x[3]&x[2]&x[1]&x[0];
assign out[3] = ~x[3]&~x[2]&~x[1]&x[0] | ~x[3]&x[2]&~x[1]&~x[0] | ~x[3]&x[2]&x[1]&x[0] |
x[3]&~x[2]&x[1]&~x[0] | x[3]&x[2]&x[1]&x[0];
assign out[4] = ~x[3]&~x[2]&~x[1]&x[0] | ~x[3]&~x[2]&x[1]&x[0] | ~x[3]&x[2]&~x[1]&~x[0] |
~x[3]&x[2]&~x[1]&x[0] | ~x[3]&x[2]&x[1]&x[0] | x[3]&~x[2]&~x[1]&x[0];
assign out[5] = ~x[3]&~x[2]&~x[1]&x[0] | ~x[3]&~x[2]&x[1]&~x[0] | ~x[3]&~x[2]&x[1]&x[0] |
~x[3]&x[2]&x[1]&x[0] | x[3]&x[2]&~x[1]&x[0];
assign out[6] = ~x[3]&~x[2]&~x[1]&~x[0] | ~x[3]&~x[2]&~x[1]&x[0] | ~x[3]&x[2]&x[1]&x[0] |
x[3]&x[2]&~x[1]&~x[0];
endmodule